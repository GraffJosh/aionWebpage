<?xml version="1.0" encoding="UTF-8"?><Batch version="2.0"><Options AppVersion="7.6.3"><PathAddFiles><![CDATA[]]></PathAddFiles><PathAddFolder><![CDATA[C:\Users\Micro\OneDrive\Projects\dev\aionWebpage\images\gallery\fullres]]></PathAddFolder></Options><TaskList><Task type="ResizeTask" enabled="true" Comment=""><Width units="1"><![CDATA[10]]></Width><Height units="1"><![CDATA[10]]></Height><DPI><![CDATA[-1]]></DPI><Filter>9</Filter><UseProportions>True</UseProportions><ResizeType>1</ResizeType><ProportionsSize>0</ProportionsSize></Task><Task type="OptimizeForWebTask" enabled="true" Comment=""><FilePath><![CDATA[C:\Users\Micro\OneDrive\Projects\dev\aionWebpage\images\gallery\previews]]></FilePath><PreserveStruct>True</PreserveStruct><CommonFolder><![CDATA[C:\Users\Micro\OneDrive\Projects\dev\aionWebpage\images\gallery\fullres\]]></CommonFolder><FileExists>1</FileExists><FileFormat>0</FileFormat><Profile>2</Profile><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGChromaSubsampling>1</JPEGChromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><JPEGRemoveMarkers>False</JPEGRemoveMarkers><JPEGProgressive>False</JPEGProgressive><JPEGBlur>0</JPEGBlur><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGTransparency>True</PNGTransparency><PNGUsePalette>False</PNGUsePalette><PNGColorCount>256</PNGColorCount><PNGInterlaced>False</PNGInterlaced><PNGRemoveTextFields>False</PNGRemoveTextFields><PNGQuality>100</PNGQuality><GIFColorCount>256</GIFColorCount><GIFTransparency>0</GIFTransparency><GIFInterlaced>0</GIFInterlaced><RemoveAllMetadata>0</RemoveAllMetadata><WEBPPreset>0</WEBPPreset><WEBPLossless>-1</WEBPLossless><WEBPQuality>100</WEBPQuality><WEBPMethod>4</WEBPMethod><WEBPTargetSize>0</WEBPTargetSize><WEBPPass>1</WEBPPass><WEBPRemoveAlpha>0</WEBPRemoveAlpha><WEBPBackColor>#FFFFFF</WEBPBackColor><WEBPAlphaQuality>100</WEBPAlphaQuality><WEBPAlphaCompression>0</WEBPAlphaCompression></Task></TaskList></Batch>